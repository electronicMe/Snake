--
--  Snake_pkg.vhd
--  The Medusa Project
--
--  Created by Sebastian Mach on 21.03.15.
--  Copyright (c) 2015. All rights reserved.
--



package Snake_pkg is

    constant numServos_c  : integer  := 26;
    constant bufferSize_c : positive := 10;

end Snake_pkg;
