--
--  Arrays_pkg.vhd
--  The Medusa Project
--
--  Created by Sebastian Mach on 06.01.15.
--  Copyright (c) 2015. All rights reserved.
--


library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;



package Arrays_pkg is

	--type NAT_ARRAY is array (integer range <>) of natural;
	type INT_ARRAY is array (integer range <>) of integer;

end;